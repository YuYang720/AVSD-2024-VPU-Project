`define CPU_CYCLE     5     // 1 Ghz
`define MAX           300000 // 30000000 cycles