`define CPU_CYCLE     1.0      // 1 Ghz
`define WDT_CYCLE     50.1     // 20 Mhz
`define MAX           30000000 // 30000000 cycles